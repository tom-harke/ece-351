stackCPU.sv